module fsm(
  input logic  [3:0] state,
  output logic [3:0] n_state
);

